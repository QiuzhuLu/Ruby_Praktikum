    1    ||  Vitello tonnato  ;  1; 15   ||   Antipasto misto   ;    1;  15   ||     Riso col nero di seppie   ;    1;  16       ||      Ossobuco ;   1;    25        ||       Panna cotta   ;   1;    7      ||   Aqua  ;  1; 10    ||       Te nero    ;    2;    4  ||     Spuma  ; 1;   4    ||     Coca    ;   1;  3    
   2  || Insalata frutti di mare    ;   1;  15     ||   Cozze al marinara  ;    1; 16  ||      Saltimboca  ;    1;    17    ||      Panna cotta ; 1;  7   ||        Tirami su  ; 1;   8     ||     Spuma   ;  2; 4     ||   Cappucino  ; 2;  4     ||     Espresso  ; 2; 4  

  3  || Antipasto misto  ;    1;   15     ||    Vitello tonnato ;    1;    15     ||     Insalata frutti di mare  ; 1;  15  ||      Saltimboca   ; 1; 17      ||   Arrosto di manzo  ;   2; 25      ||   Tirami su   ;  1;    8    ||    Caffe freddo  ;   1;    5   ||    Marsala-Zabaione  ;    1; 6     ||   Cappucino ;   2; 4     ||     Aqua   ;   2;  10       ||   Coca  ; 1;    3    



   4   ||    Insalata frutti di mare ; 2; 15        ||      Insalata mista  ;  1;    8     ||    Cozze al marinara   ;  1;    16    ||      Tirami su  ;    1;   8       ||     Coca   ;    3;   3       ||    Espresso    ;  1;  4     ||    Cappucino    ;  1;  4      ||      Spuma ;  1;  4    


    5   ||    Insalata mista    ;  1; 8   ||       Insalata frutti di mare    ;   1;   15   ||     Antipasto misto  ;   1;    15       ||      Saltimboca    ;    1;    17    ||     Cozze al marinara ;   1; 16     ||     Arrosto di manzo    ;  1;  25  ||    Tirami su   ;   1;  8   ||   Marsala-Zabaione   ;    1;   6     ||      Panna cotta   ;   1;  7        ||       Cappucino   ;    1;    4      ||    Spuma  ;    1;   4   ||    Espresso    ;   1; 4     ||   Aqua  ; 3;   10 


 6 ||    Insalata Caprese ;  2;  10   ||       Insalata frutti di mare    ; 1;   15    ||      Riso col nero di seppie  ; 1;  16    ||    Caffe freddo    ;  1;   5     ||      Marsala-Zabaione    ;    1;    6   ||     Espresso ;   3;    4       ||    Te nero ; 1;    4       ||   Coca    ;  1;   3  
  7 ||   Insalata frutti di mare ; 1;   15   ||        Cappon magro   ; 1;  28   ||       Riso col nero di seppie ;   1; 16    ||     Tirami su  ;  1;    8     ||       Marsala-Zabaione ; 1;    6    ||   Caffe freddo ; 1;    5       ||     Coca    ;  1;   3       ||   Te nero    ; 1;   4    ||   Spuma ;  1;   4 

    8  ||  Insalata frutti di mare    ;    1;    15     ||   Vitello tonnato ; 2;   15  ||    Riso col nero di seppie   ; 1; 16       ||        Pizza Margerita ;   1;   12   ||      Pizza Funghi&Salsiccia ;   1;  15       ||   Tirami su    ;  2;  8   ||       Aqua ;    3;   10      ||    Espresso   ; 1;    4    ||    Te nero   ;    1;    4    


 9  ||   Insalata frutti di mare    ; 1; 15     ||     Insalata Caprese    ;    1;    10     ||   Ossobuco    ; 1; 25  ||    Gamberoni alla griglia  ;  1; 30   ||  Panna cotta   ; 1;  7     ||       Caffe freddo    ;   1;   5    ||   Espresso  ; 1;  4     ||   Spuma ;   1;   4       ||    Te nero   ;  1; 4    

  10 || Insalata frutti di mare  ;  1;    15   ||      Antipasto misto   ;  1;  15     ||       Saltimboca ;    1;   17    ||  Pizza Margerita   ; 1;   12     ||    Caffe freddo    ;   1;    5       ||     Panna cotta   ;    1;   7   ||     Coca    ;  2;   3      ||      Te nero ;  1; 4   ||  Spuma   ;  1; 4   
